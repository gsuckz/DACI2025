** sch_path: /foss/designs/DACI2025/opamp/tb_opamp_closeloop.sch
**.subckt tb_opamp_closeloop
V1 vss GND DC{vss}
V2 vdd vss DC{vdd}
V4 vsen vcm sin(0 {vac} {fin}) dc 0 ac 1
C4 vsen vin_signal 1 m=1
I0 net1 vss DC{iref}
R1 vin vin_signal 500 m=1
R3 vout vin 5k m=1
C5 vin vss 3p m=1
C1 vout vss 20p m=1
V5 vcm vss DC{vcm}
x1 vdd net1 vin vcm vout vss v1 opamp
**** begin user architecture code




* Circuit Parameters
.param iref = 95u
.param vdd  = 1.62
.param vss  = 0.0
.param vcm  = 0.72
.param vac  = 60m
.param fin  = 9.765625e5
.options TEMP = 125.0

* FFT Parameters
.param Ts_FFT     = 1e-9
.csparam Ts_FFT   = {Ts_FFT}
.param fin_approx = 1e6
.param NFFT       = 4096
.csparam NFFT     = {NFFT}
.param vac_fin    = 'floor(fin_approx*Ts_FFT*NFFT)/Ts_FFT/NFFT'
.csparam Ti_FFT   = 3u
.csparam vac_fin  = {vac_fin}

* Include Models
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib TT
*.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red tt
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib TT
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice ss
*.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red tt
* OP Parameters & Singals to save
.save all
+ @M.X1.XM1.msky130_fd_pr__pfet_01v8_lvt[id] @M.X1.XM1.msky130_fd_pr__pfet_01v8_lvt[vth] @M.X1.XM1.msky130_fd_pr__pfet_01v8_lvt[vgs] @M.X1.XM1.msky130_fd_pr__pfet_01v8_lvt[vds] @M.X1.XM1.msky130_fd_pr__pfet_01v8_lvt[vdsat] @M.X1.XM1.msky130_fd_pr__pfet_01v8_lvt[gm] @M.X1.XM1.msky130_fd_pr__pfet_01v8_lvt[gds]
+ @M.X1.XM2.msky130_fd_pr__pfet_01v8_lvt[id] @M.X1.XM2.msky130_fd_pr__pfet_01v8_lvt[vth] @M.X1.XM2.msky130_fd_pr__pfet_01v8_lvt[vgs] @M.X1.XM2.msky130_fd_pr__pfet_01v8_lvt[vds] @M.X1.XM2.msky130_fd_pr__pfet_01v8_lvt[vdsat] @M.X1.XM2.msky130_fd_pr__pfet_01v8_lvt[gm] @M.X1.XM2.msky130_fd_pr__pfet_01v8_lvt[gds]
+ @M.X1.XM3.msky130_fd_pr__nfet_01v8[id] @M.X1.XM3.msky130_fd_pr__nfet_01v8[vth] @M.X1.XM3.msky130_fd_pr__nfet_01v8[vgs] @M.X1.XM3.msky130_fd_pr__nfet_01v8[vds] @M.X1.XM3.msky130_fd_pr__nfet_01v8[vdsat] @M.X1.XM3.msky130_fd_pr__nfet_01v8[gm] @M.X1.XM3.msky130_fd_pr__nfet_01v8[gds]
+ @M.X1.XM4.msky130_fd_pr__nfet_01v8[id] @M.X1.XM4.msky130_fd_pr__nfet_01v8[vth] @M.X1.XM4.msky130_fd_pr__nfet_01v8[vgs] @M.X1.XM4.msky130_fd_pr__nfet_01v8[vds] @M.X1.XM4.msky130_fd_pr__nfet_01v8[vdsat] @M.X1.XM4.msky130_fd_pr__nfet_01v8[gm] @M.X1.XM4.msky130_fd_pr__nfet_01v8[gds]
+ @M.X1.XM5.msky130_fd_pr__pfet_01v8[id] @M.X1.XM5.msky130_fd_pr__pfet_01v8[vth] @M.X1.XM5.msky130_fd_pr__pfet_01v8[vgs] @M.X1.XM5.msky130_fd_pr__pfet_01v8[vds] @M.X1.XM5.msky130_fd_pr__pfet_01v8[vdsat] @M.X1.XM5.msky130_fd_pr__pfet_01v8[gm] @M.X1.XM5.msky130_fd_pr__pfet_01v8[gds]
+ @M.X1.XM6.msky130_fd_pr__nfet_01v8[id] @M.X1.XM6.msky130_fd_pr__nfet_01v8[vth] @M.X1.XM6.msky130_fd_pr__nfet_01v8[vgs] @M.X1.XM6.msky130_fd_pr__nfet_01v8[vds] @M.X1.XM6.msky130_fd_pr__nfet_01v8[vdsat] @M.X1.XM6.msky130_fd_pr__nfet_01v8[gm] @M.X1.XM6.msky130_fd_pr__nfet_01v8[gds]
+ @M.X1.XM7.msky130_fd_pr__pfet_01v8[id] @M.X1.XM7.msky130_fd_pr__pfet_01v8[vth] @M.X1.XM7.msky130_fd_pr__pfet_01v8[vgs] @M.X1.XM7.msky130_fd_pr__pfet_01v8[vds] @M.X1.XM7.msky130_fd_pr__pfet_01v8[vdsat] @M.X1.XM7.msky130_fd_pr__pfet_01v8[gm] @M.X1.XM7.msky130_fd_pr__pfet_01v8[gds]
+ @M.X1.XM8.msky130_fd_pr__pfet_01v8[id] @M.X1.XM8.msky130_fd_pr__pfet_01v8[vth] @M.X1.XM8.msky130_fd_pr__pfet_01v8[vgs] @M.X1.XM8.msky130_fd_pr__pfet_01v8[vds] @M.X1.XM8.msky130_fd_pr__pfet_01v8[vdsat] @M.X1.XM8.msky130_fd_pr__pfet_01v8[gm] @M.X1.XM8.msky130_fd_pr__pfet_01v8[gds]
+ @M.X1.XM9.msky130_fd_pr__nfet_01v8[id] @M.X1.XM9.msky130_fd_pr__nfet_01v8[vth] @M.X1.XM9.msky130_fd_pr__nfet_01v8[vgs] @M.X1.XM9.msky130_fd_pr__nfet_01v8[vds] @M.X1.XM9.msky130_fd_pr__nfet_01v8[vdsat] @M.X1.XM9.msky130_fd_pr__nfet_01v8[gm] @M.X1.XM9.msky130_fd_pr__nfet_01v8[gds]

*Simulation
.control
  set color0 = white

  ac dec 100 1k 10G
  setplot ac1
  meas ac GBW when vdb(vout)=0
  meas ac DCG find vdb(vout) at=1k
  meas ac PM find vp(vout) when vdb(vout)=0
  print PM*180/PI
  plot vdb(vout) {vp(vout)*180/PI} vdb(v1) {vp(v1)*180/PI}

  reset
  tran 0.01u 11u
  setplot tran1
  plot v(vsen) v(vout)

  *reset
  *set sqrnoise
  *noise v(vout) V4 dec 100 1k 10G 1
  *let onoise_total_integrado = maximum(sqrt(integ(onoise_spectrum)))
  *print onoise_total_integrado



  reset
  tran 0.001u 11u
  fourier 9.765625e5 vout
  let THD_db = db(fourier11[1][3]/fourier11[1][1])
  print THD_db
  let lin-tstart = {Ti_FFT} $ skip the start - up phase
  let lin-tstep = {Ts_FFT}
  let lin-tstop = {Ti_FFT + (NFFT-1) * Ts_FFT} $ end earlier
  linearize vout
  set specwindow = none
 fft vout
  plot mag(vout)
  plot db(mag(vout)) xlimit 0 20e6

  reset
  op
  setplot op1
  unset filetype
  write tb_opamp_closeloop.raw


  reset
  noise v(vout) V4 dec 100 1k 10G 1
  setplot noise1
  plot onoise_spectrum
  setplot noise2
  print inoise_total
  print onoise_total
  print onoise_total.m.x1.xm1.msky130_fd_pr__pfet_01v8_lvt.1overf
  print onoise_total.m.x1.xm1.msky130_fd_pr__pfet_01v8_lvt.id
  print onoise_total.m.x1.xm2.msky130_fd_pr__pfet_01v8_lvt.1overf
  print onoise_total.m.x1.xm2.msky130_fd_pr__pfet_01v8_lvt.id
  print onoise_total.m.x1.xm3.msky130_fd_pr__nfet_01v8.1overf
  print onoise_total.m.x1.xm3.msky130_fd_pr__nfet_01v8.id
  print onoise_total.m.x1.xm4.msky130_fd_pr__nfet_01v8.1overf
  print onoise_total.m.x1.xm4.msky130_fd_pr__nfet_01v8.id
  print onoise_total.m.x1.xm5.msky130_fd_pr__pfet_01v8.1overf
  print onoise_total.m.x1.xm5.msky130_fd_pr__pfet_01v8.id
  print onoise_total.m.x1.xm6.msky130_fd_pr__nfet_01v8.1overf
  print onoise_total.m.x1.xm6.msky130_fd_pr__nfet_01v8.id
  print onoise_total.m.x1.xm7.msky130_fd_pr__pfet_01v8.1overf
  print onoise_total.m.x1.xm7.msky130_fd_pr__pfet_01v8.id
  vprint onoise_total.m.x1.xm8.msky130_fd_pr__pfet_01v8.1overf
  print onoise_total.m.x1.xm8.msky130_fd_pr__pfet_01v8.id
  set filetype=ascii
  write tpfinal_noise.raw
.endc

.end


**** end user architecture code
**.ends

* expanding   symbol:  opamp.sym # of pins=7
** sym_path: /foss/designs/DACI2025/opamp/opamp.sym
** sch_path: /foss/designs/DACI2025/opamp/opamp.sch
.subckt opamp vdd iref vin_n vin_p vout vss v1
*.iopin vdd
*.iopin vss
*.ipin vin_n
*.ipin vin_p
*.ipin iref
*.opin vout
*.opin v1
XM5 vp iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=50 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=27 m=27
XM7 vout iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=50 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24
XM8 iref iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=50 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
XM1 vbn vin_n vp vp sky130_fd_pr__pfet_01v8_lvt L=0.6 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM2 v1 vin_p vp vp sky130_fd_pr__pfet_01v8_lvt L=0.6 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
C1 net2 vout 7.9p m=1
Vmeas net1 vss 0
.save i(vmeas)
R7 net2 v1 350 m=1
XM6 vout v1 net1 net1 sky130_fd_pr__nfet_01v8 L=0.3 W=35 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM4 v1 vbn net1 net1 sky130_fd_pr__nfet_01v8 L=2.2 W=80 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 vbn vbn net1 net1 sky130_fd_pr__nfet_01v8 L=2.2 W=80 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends

.GLOBAL GND
.end
