** sch_path: /foss/designs/DACI2025/tp3/tp3_1.sch
**.subckt tp3_1
Iref vdd vbn {iref}
VSS vss GND {vss}
VDD vdd vss {vdd}
V1 net1 vss {vcm}
XM1 net2 vbn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.75 W={wn} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM0 vbn vbn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.75 W={wn} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM2 vout1 vin1 net2 vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W={wdif} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R2 vdd vout1 {R} m=1
XM3 vout2 vin2 net2 vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W={wdif} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R1 vdd vout2 {R} m=1
V2 vin1 net1 SIN(0 {Vin} 50Meg) DC 0
V3 net1 vin2 SIN(0 {Vin} 50Meg) DC 0 AC 1
**** begin user architecture code



* Parameters
.param vdd = 1.8
.param vss = 0.0
.param iref = 100u
.param wn = 8
.param wdif = 3.5
.param R = 12k
.param Vin = 10m
.param vcm = 1.2

.options TEMP = 65.0

* Models
*.lib ~/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/sky130.lib TT
*.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red tt
* Data to save
.save all
+ @M.XM0.msky130_fd_pr__nfet_01v8_lvt[id]
+ @M.XM0.msky130_fd_pr__nfet_01v8_lvt[vds]
+ @M.XM0.msky130_fd_pr__nfet_01v8_lvt[vgs]
+ @M.XM0.msky130_fd_pr__nfet_01v8_lvt[vdsat]
+ @M.XM0.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @M.XM0.msky130_fd_pr__nfet_01v8_lvt[gm]
+ @M.XM1.msky130_fd_pr__nfet_01v8_lvt[id]
+ @M.XM1.msky130_fd_pr__nfet_01v8_lvt[vds]
+ @M.XM1.msky130_fd_pr__nfet_01v8_lvt[vgs]
+ @M.XM1.msky130_fd_pr__nfet_01v8_lvt[vdsat]
+ @M.XM1.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @M.XM1.msky130_fd_pr__nfet_01v8_lvt[gm]
+ @M.XM1.msky130_fd_pr__nfet_01v8_lvt[gds]
+ @M.XM2.msky130_fd_pr__nfet_01v8_lvt[id]
+ @M.XM2.msky130_fd_pr__nfet_01v8_lvt[vds]
+ @M.XM2.msky130_fd_pr__nfet_01v8_lvt[vgs]
+ @M.XM2.msky130_fd_pr__nfet_01v8_lvt[vdsat]
+ @M.XM2.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @M.XM2.msky130_fd_pr__nfet_01v8_lvt[gm]
+ @M.XM2.msky130_fd_pr__nfet_01v8_lvt[gds]
+ @M.XM3.msky130_fd_pr__nfet_01v8_lvt[id]
+ @M.XM3.msky130_fd_pr__nfet_01v8_lvt[vds]
+ @M.XM3.msky130_fd_pr__nfet_01v8_lvt[vgs]
+ @M.XM3.msky130_fd_pr__nfet_01v8_lvt[vdsat]
+ @M.XM3.msky130_fd_pr__nfet_01v8_lvt[vth]
+ @M.XM3.msky130_fd_pr__nfet_01v8_lvt[gm]
+ @M.XM3.msky130_fd_pr__nfet_01v8_lvt[gds]

* Simulation
.control


  ac dec 100 10k 100G
  let vdiff = vout1-vout2
  let vindiff = vin1-vin2
  setplot ac1
  meas ac GBW when vdb(vdiff) = 0
  meas ac DCG find vdb(vdiff) at=10k
  meas ac PM find vp(vdiff) when vdb(vdiff)=0
  print PM*180/PI
  meas ac GM find vdb(vdiff) when vp(vdiff)=0
  plot vdb(vdiff) {vp(vdiff)*180/PI}
  write tp3_1_ac.raw

  reset
  tran 0.01n 100n
  let vdiff = vout1-vout2
  let vindiff = vin1-vin2
  plot v(vindiff) v(vdiff)
 plot v(vout1) v(vout2)
 plot v(vin1) v(vin2)
  write tp3_1_tran.raw
reset
 op
  save all
  print all
  unset filetype
  write tp3_1.raw



.endc

.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
