** sch_path: /foss/designs/DACI2025/opamp/untitled.sch
**.subckt untitled
**.ends
.end
